`default_nettype none
`timescale 1ns / 1ps

module eth_packer (
    input wire clk,
    input wire rst,
    input wire axiiv,
    input wire [7:0] pixel,

    output logic phy_txen,
    output logic [1:0] phy_txd
);
logic [3:0] state;
logic [2:0] byte_bit_counter;
logic [12:0] dibit_counter;

always_comb begin
    if (axiiv) begin

    end
end

always_ff(@posedge clk) begin

end


endmodule

`default_nettype wire